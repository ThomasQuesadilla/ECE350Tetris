`define VIDEO_WIDTH 640  // Standard VGA Width
`define VIDEO_HEIGHT 480 // Standard VGA Height

`define PLAYAREA_START 200
`define PLAYAREA_END 440